module spi_master (

);

endmodule