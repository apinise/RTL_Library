module i2c_slave (

);

endmodule