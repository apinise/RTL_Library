module mux_hot #(
  parameter INPUTS  = 2,
  parameter WIDTH   = 32
)(
  input   logic [WIDTH-1:0]   inputs [INPUTS],
  input   logic [INPUTS-1:0]  sel,
  output  logic [WIDTH-1:0]   out
);

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

integer i;

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

always_comb begin
  out = 'z;
  for (i=0; i<INPUTS; i=i+1) begin
    if (sel == (1 << i)) begin
      out = inputs[i];
    end
  end
end

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////
/*
mux_hot mux #(
  .INPUTS(),
  .WIDTH()
)(
  .inputs(),
  .sel(),
  .out()
);
*/

endmodule